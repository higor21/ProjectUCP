library verilog;
use verilog.vl_types.all;
entity Processador_vlg_check_tst is
    port(
        Q1              : in     vl_logic_vector(6 downto 0);
        Q2              : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end Processador_vlg_check_tst;
